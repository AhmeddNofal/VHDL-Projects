--
-- VHDL Architecture my_project_lib.encoder.rtl
--
-- Created:
--          by - Owner.UNKNOWN (DESKTOP-BED4071)
--          at - 17:43:21 12/ 2/2022
--
-- using Mentor Graphics HDL Designer(TM) 2007.1 (Build 19)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY encoder IS
  port ( a : in std_logic_vector(7 downto 0);
         y : out std_logic_vector(2 downto 0));
END ENTITY encoder;

--
ARCHITECTURE rtl OF encoder IS
BEGIN
  with a select 
    y<= "000" when "00000001",
        "001" when "00000010",
        "010" when "00000100",
        "011" when "00001000",
        "100" when "00010000",
        "101" when "00100000",
        "110" when "01000000",
        "111" when "10000000",
        "---" when others;
END ARCHITECTURE rtl;

